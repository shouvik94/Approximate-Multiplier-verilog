module test;
    reg[7:0] a,b;
    wire[10:0] out;

    main_mul m1(a,b,out);
    initial begin
        #5 a=8'b01011011;b=8'b01110101;
        #5 a=8'b00000001;b=8'b00000001;
        #5 a=8'b11111111;b=8'b11111111;
        #5 a=8'b01001000;b=8'b11100101;
        #5 a=8'b10010111;b=8'b10000010;
        #5 a=8'b11110101;b=8'b00011111;
        #5 a=8'b01010101;b=8'b01111110;
        #5 a=8'b00110101;b=8'b00000000;
        #5 a=8'b01011111;b=8'b00111100;
        #5 a=8'b11010110;b=8'b11001010;
        #5 a=8'b01111111;b=8'b01111111;
    end
    
    always @(out)
    begin
        $display("A=%b,B=%b,Out=%b",a,b,out);
    end

endmodule